
-- In this example, we're going to map voltage to distance, using a linear 
-- approximation, according to the Sharp GP2Y0A41SK0F datasheet page 4, or 
-- Lab 3 handout page 5. 
-- 
-- The relevant points we will select are:
-- 2.750 V is  4.00 cm (or 2750 mV and  40.0 mm)
-- 0.400 V is 33.00 cm (or  400 mV and 330.0 mm)
-- 
-- Mapping to the scales in our system
-- 2750 (mV) should map to  400 (10^-4 m)
--  400 (mV) should map to 3300 (10^-4 m)
-- and developing a linear equation, we find:
--
-- Distance = -2900/2350 * Voltage + 3793.617
-- Note this code implements linear function, you must map to the 
-- NON-linear relationship in the datasheet. This code is only provided 
-- for reference to help get you started.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY voltage2distance IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      voltage        :  IN    STD_LOGIC_VECTOR(12 DOWNTO 0);                           
      distance       :  OUT   STD_LOGIC_VECTOR(12 DOWNTO 0));  
END voltage2distance;

ARCHITECTURE behavior OF voltage2distance IS

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.
-- See how to get the distance output at the bottom of this file,
-- after begin.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3333	)	,
(	3297	)	,
(	3290	)	,
(	3282	)	,
(	3275	)	,
(	3268	)	,
(	3260	)	,
(	3253	)	,
(	3246	)	,
(	3239	)	,
(	3232	)	,
(	3225	)	,
(	3218	)	,
(	3211	)	,
(	3203	)	,
(	3196	)	,
(	3189	)	,
(	3182	)	,
(	3175	)	,
(	3169	)	,
(	3162	)	,
(	3155	)	,
(	3148	)	,
(	3141	)	,
(	3134	)	,
(	3127	)	,
(	3121	)	,
(	3114	)	,
(	3107	)	,
(	3100	)	,
(	3094	)	,
(	3087	)	,
(	3080	)	,
(	3074	)	,
(	3067	)	,
(	3060	)	,
(	3054	)	,
(	3047	)	,
(	3041	)	,
(	3034	)	,
(	3028	)	,
(	3021	)	,
(	3015	)	,
(	3008	)	,
(	3002	)	,
(	2996	)	,
(	2989	)	,
(	2983	)	,
(	2977	)	,
(	2970	)	,
(	2964	)	,
(	2958	)	,
(	2951	)	,
(	2945	)	,
(	2939	)	,
(	2933	)	,
(	2927	)	,
(	2920	)	,
(	2914	)	,
(	2908	)	,
(	2902	)	,
(	2896	)	,
(	2890	)	,
(	2884	)	,
(	2878	)	,
(	2872	)	,
(	2866	)	,
(	2860	)	,
(	2854	)	,
(	2848	)	,
(	2842	)	,
(	2836	)	,
(	2830	)	,
(	2825	)	,
(	2819	)	,
(	2813	)	,
(	2807	)	,
(	2801	)	,
(	2796	)	,
(	2790	)	,
(	2784	)	,
(	2778	)	,
(	2773	)	,
(	2767	)	,
(	2761	)	,
(	2756	)	,
(	2750	)	,
(	2745	)	,
(	2739	)	,
(	2733	)	,
(	2728	)	,
(	2722	)	,
(	2717	)	,
(	2711	)	,
(	2706	)	,
(	2700	)	,
(	2695	)	,
(	2689	)	,
(	2684	)	,
(	2679	)	,
(	2673	)	,
(	2668	)	,
(	2663	)	,
(	2657	)	,
(	2652	)	,
(	2647	)	,
(	2641	)	,
(	2636	)	,
(	2631	)	,
(	2626	)	,
(	2620	)	,
(	2615	)	,
(	2610	)	,
(	2605	)	,
(	2600	)	,
(	2595	)	,
(	2590	)	,
(	2585	)	,
(	2579	)	,
(	2574	)	,
(	2569	)	,
(	2564	)	,
(	2559	)	,
(	2554	)	,
(	2549	)	,
(	2544	)	,
(	2539	)	,
(	2534	)	,
(	2530	)	,
(	2525	)	,
(	2520	)	,
(	2515	)	,
(	2510	)	,
(	2505	)	,
(	2500	)	,
(	2496	)	,
(	2491	)	,
(	2486	)	,
(	2481	)	,
(	2476	)	,
(	2472	)	,
(	2467	)	,
(	2462	)	,
(	2458	)	,
(	2453	)	,
(	2448	)	,
(	2444	)	,
(	2439	)	,
(	2434	)	,
(	2430	)	,
(	2425	)	,
(	2421	)	,
(	2416	)	,
(	2411	)	,
(	2407	)	,
(	2402	)	,
(	2398	)	,
(	2393	)	,
(	2389	)	,
(	2385	)	,
(	2380	)	,
(	2376	)	,
(	2371	)	,
(	2367	)	,
(	2362	)	,
(	2358	)	,
(	2354	)	,
(	2349	)	,
(	2345	)	,
(	2341	)	,
(	2336	)	,
(	2332	)	,
(	2328	)	,
(	2324	)	,
(	2319	)	,
(	2315	)	,
(	2311	)	,
(	2307	)	,
(	2302	)	,
(	2298	)	,
(	2294	)	,
(	2290	)	,
(	2286	)	,
(	2282	)	,
(	2277	)	,
(	2273	)	,
(	2269	)	,
(	2265	)	,
(	2261	)	,
(	2257	)	,
(	2253	)	,
(	2249	)	,
(	2245	)	,
(	2241	)	,
(	2237	)	,
(	2233	)	,
(	2229	)	,
(	2225	)	,
(	2221	)	,
(	2217	)	,
(	2213	)	,
(	2209	)	,
(	2205	)	,
(	2202	)	,
(	2198	)	,
(	2194	)	,
(	2190	)	,
(	2186	)	,
(	2182	)	,
(	2179	)	,
(	2175	)	,
(	2171	)	,
(	2167	)	,
(	2163	)	,
(	2160	)	,
(	2156	)	,
(	2152	)	,
(	2148	)	,
(	2145	)	,
(	2141	)	,
(	2137	)	,
(	2134	)	,
(	2130	)	,
(	2126	)	,
(	2123	)	,
(	2119	)	,
(	2115	)	,
(	2112	)	,
(	2108	)	,
(	2105	)	,
(	2101	)	,
(	2098	)	,
(	2094	)	,
(	2090	)	,
(	2087	)	,
(	2083	)	,
(	2080	)	,
(	2076	)	,
(	2073	)	,
(	2069	)	,
(	2066	)	,
(	2063	)	,
(	2059	)	,
(	2056	)	,
(	2052	)	,
(	2049	)	,
(	2045	)	,
(	2042	)	,
(	2039	)	,
(	2035	)	,
(	2032	)	,
(	2029	)	,
(	2025	)	,
(	2022	)	,
(	2019	)	,
(	2015	)	,
(	2012	)	,
(	2009	)	,
(	2006	)	,
(	2002	)	,
(	1999	)	,
(	1996	)	,
(	1993	)	,
(	1989	)	,
(	1986	)	,
(	1983	)	,
(	1980	)	,
(	1976	)	,
(	1973	)	,
(	1970	)	,
(	1967	)	,
(	1964	)	,
(	1961	)	,
(	1958	)	,
(	1954	)	,
(	1951	)	,
(	1948	)	,
(	1945	)	,
(	1942	)	,
(	1939	)	,
(	1936	)	,
(	1933	)	,
(	1930	)	,
(	1927	)	,
(	1924	)	,
(	1921	)	,
(	1918	)	,
(	1915	)	,
(	1912	)	,
(	1909	)	,
(	1906	)	,
(	1903	)	,
(	1900	)	,
(	1897	)	,
(	1894	)	,
(	1891	)	,
(	1888	)	,
(	1885	)	,
(	1882	)	,
(	1879	)	,
(	1877	)	,
(	1874	)	,
(	1871	)	,
(	1868	)	,
(	1865	)	,
(	1862	)	,
(	1859	)	,
(	1857	)	,
(	1854	)	,
(	1851	)	,
(	1848	)	,
(	1845	)	,
(	1843	)	,
(	1840	)	,
(	1837	)	,
(	1834	)	,
(	1832	)	,
(	1829	)	,
(	1826	)	,
(	1823	)	,
(	1821	)	,
(	1818	)	,
(	1815	)	,
(	1813	)	,
(	1810	)	,
(	1807	)	,
(	1805	)	,
(	1802	)	,
(	1799	)	,
(	1797	)	,
(	1794	)	,
(	1791	)	,
(	1789	)	,
(	1786	)	,
(	1783	)	,
(	1781	)	,
(	1778	)	,
(	1776	)	,
(	1773	)	,
(	1771	)	,
(	1768	)	,
(	1765	)	,
(	1763	)	,
(	1760	)	,
(	1758	)	,
(	1755	)	,
(	1753	)	,
(	1750	)	,
(	1748	)	,
(	1745	)	,
(	1743	)	,
(	1740	)	,
(	1738	)	,
(	1735	)	,
(	1733	)	,
(	1730	)	,
(	1728	)	,
(	1726	)	,
(	1723	)	,
(	1721	)	,
(	1718	)	,
(	1716	)	,
(	1713	)	,
(	1711	)	,
(	1709	)	,
(	1706	)	,
(	1704	)	,
(	1702	)	,
(	1699	)	,
(	1697	)	,
(	1695	)	,
(	1692	)	,
(	1690	)	,
(	1688	)	,
(	1685	)	,
(	1683	)	,
(	1681	)	,
(	1678	)	,
(	1676	)	,
(	1674	)	,
(	1671	)	,
(	1669	)	,
(	1667	)	,
(	1665	)	,
(	1662	)	,
(	1660	)	,
(	1658	)	,
(	1656	)	,
(	1653	)	,
(	1651	)	,
(	1649	)	,
(	1647	)	,
(	1644	)	,
(	1642	)	,
(	1640	)	,
(	1638	)	,
(	1636	)	,
(	1634	)	,
(	1631	)	,
(	1629	)	,
(	1627	)	,
(	1625	)	,
(	1623	)	,
(	1621	)	,
(	1618	)	,
(	1616	)	,
(	1614	)	,
(	1612	)	,
(	1610	)	,
(	1608	)	,
(	1606	)	,
(	1604	)	,
(	1602	)	,
(	1599	)	,
(	1597	)	,
(	1595	)	,
(	1593	)	,
(	1591	)	,
(	1589	)	,
(	1587	)	,
(	1585	)	,
(	1583	)	,
(	1581	)	,
(	1579	)	,
(	1577	)	,
(	1575	)	,
(	1573	)	,
(	1571	)	,
(	1569	)	,
(	1567	)	,
(	1565	)	,
(	1563	)	,
(	1561	)	,
(	1559	)	,
(	1557	)	,
(	1555	)	,
(	1553	)	,
(	1551	)	,
(	1549	)	,
(	1547	)	,
(	1545	)	,
(	1543	)	,
(	1541	)	,
(	1540	)	,
(	1538	)	,
(	1536	)	,
(	1534	)	,
(	1532	)	,
(	1530	)	,
(	1528	)	,
(	1526	)	,
(	1524	)	,
(	1522	)	,
(	1521	)	,
(	1519	)	,
(	1517	)	,
(	1515	)	,
(	1513	)	,
(	1511	)	,
(	1509	)	,
(	1508	)	,
(	1506	)	,
(	1504	)	,
(	1502	)	,
(	1500	)	,
(	1498	)	,
(	1497	)	,
(	1495	)	,
(	1493	)	,
(	1491	)	,
(	1489	)	,
(	1488	)	,
(	1486	)	,
(	1484	)	,
(	1482	)	,
(	1481	)	,
(	1479	)	,
(	1477	)	,
(	1475	)	,
(	1473	)	,
(	1472	)	,
(	1470	)	,
(	1468	)	,
(	1466	)	,
(	1465	)	,
(	1463	)	,
(	1461	)	,
(	1460	)	,
(	1458	)	,
(	1456	)	,
(	1454	)	,
(	1453	)	,
(	1451	)	,
(	1449	)	,
(	1448	)	,
(	1446	)	,
(	1444	)	,
(	1443	)	,
(	1441	)	,
(	1439	)	,
(	1438	)	,
(	1436	)	,
(	1434	)	,
(	1433	)	,
(	1431	)	,
(	1429	)	,
(	1428	)	,
(	1426	)	,
(	1424	)	,
(	1423	)	,
(	1421	)	,
(	1420	)	,
(	1418	)	,
(	1416	)	,
(	1415	)	,
(	1413	)	,
(	1412	)	,
(	1410	)	,
(	1408	)	,
(	1407	)	,
(	1405	)	,
(	1404	)	,
(	1402	)	,
(	1400	)	,
(	1399	)	,
(	1397	)	,
(	1396	)	,
(	1394	)	,
(	1393	)	,
(	1391	)	,
(	1389	)	,
(	1388	)	,
(	1386	)	,
(	1385	)	,
(	1383	)	,
(	1382	)	,
(	1380	)	,
(	1379	)	,
(	1377	)	,
(	1376	)	,
(	1374	)	,
(	1373	)	,
(	1371	)	,
(	1370	)	,
(	1368	)	,
(	1367	)	,
(	1365	)	,
(	1364	)	,
(	1362	)	,
(	1361	)	,
(	1359	)	,
(	1358	)	,
(	1356	)	,
(	1355	)	,
(	1353	)	,
(	1352	)	,
(	1350	)	,
(	1349	)	,
(	1347	)	,
(	1346	)	,
(	1345	)	,
(	1343	)	,
(	1342	)	,
(	1340	)	,
(	1339	)	,
(	1337	)	,
(	1336	)	,
(	1334	)	,
(	1333	)	,
(	1332	)	,
(	1330	)	,
(	1329	)	,
(	1327	)	,
(	1326	)	,
(	1325	)	,
(	1323	)	,
(	1322	)	,
(	1320	)	,
(	1319	)	,
(	1318	)	,
(	1316	)	,
(	1315	)	,
(	1313	)	,
(	1312	)	,
(	1311	)	,
(	1309	)	,
(	1308	)	,
(	1307	)	,
(	1305	)	,
(	1304	)	,
(	1302	)	,
(	1301	)	,
(	1300	)	,
(	1298	)	,
(	1297	)	,
(	1296	)	,
(	1294	)	,
(	1293	)	,
(	1292	)	,
(	1290	)	,
(	1289	)	,
(	1288	)	,
(	1286	)	,
(	1285	)	,
(	1284	)	,
(	1282	)	,
(	1281	)	,
(	1280	)	,
(	1278	)	,
(	1277	)	,
(	1276	)	,
(	1274	)	,
(	1273	)	,
(	1272	)	,
(	1271	)	,
(	1269	)	,
(	1268	)	,
(	1267	)	,
(	1265	)	,
(	1264	)	,
(	1263	)	,
(	1262	)	,
(	1260	)	,
(	1259	)	,
(	1258	)	,
(	1256	)	,
(	1255	)	,
(	1254	)	,
(	1253	)	,
(	1251	)	,
(	1250	)	,
(	1249	)	,
(	1248	)	,
(	1246	)	,
(	1245	)	,
(	1244	)	,
(	1243	)	,
(	1241	)	,
(	1240	)	,
(	1239	)	,
(	1238	)	,
(	1237	)	,
(	1235	)	,
(	1234	)	,
(	1233	)	,
(	1232	)	,
(	1230	)	,
(	1229	)	,
(	1228	)	,
(	1227	)	,
(	1226	)	,
(	1224	)	,
(	1223	)	,
(	1222	)	,
(	1221	)	,
(	1220	)	,
(	1218	)	,
(	1217	)	,
(	1216	)	,
(	1215	)	,
(	1214	)	,
(	1212	)	,
(	1211	)	,
(	1210	)	,
(	1209	)	,
(	1208	)	,
(	1206	)	,
(	1205	)	,
(	1204	)	,
(	1203	)	,
(	1202	)	,
(	1201	)	,
(	1199	)	,
(	1198	)	,
(	1197	)	,
(	1196	)	,
(	1195	)	,
(	1194	)	,
(	1193	)	,
(	1191	)	,
(	1190	)	,
(	1189	)	,
(	1188	)	,
(	1187	)	,
(	1186	)	,
(	1185	)	,
(	1183	)	,
(	1182	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1178	)	,
(	1177	)	,
(	1175	)	,
(	1174	)	,
(	1173	)	,
(	1172	)	,
(	1171	)	,
(	1170	)	,
(	1169	)	,
(	1168	)	,
(	1167	)	,
(	1165	)	,
(	1164	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1159	)	,
(	1158	)	,
(	1157	)	,
(	1156	)	,
(	1155	)	,
(	1153	)	,
(	1152	)	,
(	1151	)	,
(	1150	)	,
(	1149	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1145	)	,
(	1144	)	,
(	1143	)	,
(	1142	)	,
(	1141	)	,
(	1140	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1134	)	,
(	1133	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1127	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1121	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1114	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1099	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1090	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1025	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1010	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	991	)	,
(	990	)	,
(	989	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	985	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	976	)	,
(	975	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	972	)	,
(	971	)	,
(	970	)	,
(	970	)	,
(	969	)	,
(	968	)	,
(	967	)	,
(	966	)	,
(	966	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	962	)	,
(	961	)	,
(	961	)	,
(	960	)	,
(	959	)	,
(	958	)	,
(	957	)	,
(	957	)	,
(	956	)	,
(	955	)	,
(	954	)	,
(	953	)	,
(	953	)	,
(	952	)	,
(	951	)	,
(	950	)	,
(	949	)	,
(	949	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	945	)	,
(	945	)	,
(	944	)	,
(	943	)	,
(	942	)	,
(	941	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	938	)	,
(	938	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	934	)	,
(	934	)	,
(	933	)	,
(	932	)	,
(	931	)	,
(	931	)	,
(	930	)	,
(	929	)	,
(	928	)	,
(	927	)	,
(	927	)	,
(	926	)	,
(	925	)	,
(	924	)	,
(	924	)	,
(	923	)	,
(	922	)	,
(	921	)	,
(	921	)	,
(	920	)	,
(	919	)	,
(	918	)	,
(	918	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	915	)	,
(	914	)	,
(	913	)	,
(	912	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	909	)	,
(	909	)	,
(	908	)	,
(	907	)	,
(	906	)	,
(	906	)	,
(	905	)	,
(	904	)	,
(	903	)	,
(	903	)	,
(	902	)	,
(	901	)	,
(	900	)	,
(	900	)	,
(	899	)	,
(	898	)	,
(	897	)	,
(	897	)	,
(	896	)	,
(	895	)	,
(	895	)	,
(	894	)	,
(	893	)	,
(	892	)	,
(	892	)	,
(	891	)	,
(	890	)	,
(	889	)	,
(	889	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	885	)	,
(	884	)	,
(	884	)	,
(	883	)	,
(	882	)	,
(	882	)	,
(	881	)	,
(	880	)	,
(	879	)	,
(	879	)	,
(	878	)	,
(	877	)	,
(	877	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	868	)	,
(	867	)	,
(	866	)	,
(	866	)	,
(	865	)	,
(	864	)	,
(	863	)	,
(	863	)	,
(	862	)	,
(	861	)	,
(	861	)	,
(	860	)	,
(	859	)	,
(	859	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	855	)	,
(	855	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	851	)	,
(	851	)	,
(	850	)	,
(	849	)	,
(	849	)	,
(	848	)	,
(	847	)	,
(	847	)	,
(	846	)	,
(	845	)	,
(	845	)	,
(	844	)	,
(	843	)	,
(	843	)	,
(	842	)	,
(	841	)	,
(	841	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	837	)	,
(	837	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	834	)	,
(	833	)	,
(	832	)	,
(	832	)	,
(	831	)	,
(	830	)	,
(	830	)	,
(	829	)	,
(	828	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	823	)	,
(	823	)	,
(	822	)	,
(	821	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	815	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	812	)	,
(	811	)	,
(	810	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	804	)	,
(	803	)	,
(	802	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	797	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	794	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	785	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	755	)	,
(	754	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	742	)	,
(	741	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	713	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	705	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	702	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	696	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	684	)	,
(	683	)	,
(	683	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	681	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	676	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	672	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	669	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	658	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	654	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	639	)	,
(	639	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	637	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	635	)	,
(	635	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	633	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	629	)	,
(	629	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	626	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	622	)	,
(	622	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	619	)	,
(	619	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	617	)	,
(	617	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	613	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	610	)	,
(	610	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	607	)	,
(	607	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	601	)	,
(	601	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	596	)	,
(	596	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	592	)	,
(	592	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	589	)	,
(	589	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	586	)	,
(	586	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	582	)	,
(	582	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	579	)	,
(	579	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	570	)	,
(	570	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	564	)	,
(	564	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	559	)	,
(	559	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	


);


begin
   -- This is the only statement required. It looks up the converted value of 
	-- the voltage input (in mV) in the v2d_LUT look-up table, and outputs the 
	-- distance (in 10^-4 m) in std_logic_vector format.
    	
   distance <= std_logic_vector(to_unsigned(v2d_LUT(to_integer(unsigned(voltage))),distance'length));

end behavior;